// megafunction wizard: %ALTPLL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altpll

// ============================================================
// File Name: pll.v
// Megafunction Name(s):
// 			altpll
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module pll (
           inclk0,
           c0);

input	  inclk0;
output	  c0;

wire [5:0] sub_wire0;
wire [0:0] sub_wire4 = 1'h0;
wire [0:0] sub_wire1 = sub_wire0[0:0];
wire  c0 = sub_wire1;
wire  sub_wire2 = inclk0;
wire [1:0] sub_wire3 = {sub_wire4, sub_wire2};

altpll	altpll_component (
           .inclk (sub_wire3),
           .clk (sub_wire0),
           .activeclock (),
           .areset (1'b0),
           .clkbad (),
           .clkena ({6{1'b1}}),
           .clkloss (),
           .clkswitch (1'b0),
           .configupdate (1'b0),
           .enable0 (),
           .enable1 (),
           .extclk (),
           .extclkena ({4{1'b1}}),
           .fbin (1'b1),
           .fbmimicbidir (),
           .fbout (),
           .fref (),
           .icdrclk (),
           .locked (),
           .pfdena (1'b1),
           .phasecounterselect ({4{1'b1}}),
           .phasedone (),
           .phasestep (1'b1),
           .phaseupdown (1'b1),
           .pllena (1'b1),
           .scanaclr (1'b0),
           .scanclk (1'b0),
           .scanclkena (1'b1),
           .scandata (1'b0),
           .scandataout (),
           .scandone (),
           .scanread (1'b0),
           .scanwrite (1'b0),
           .sclkout0 (),
           .sclkout1 (),
           .vcooverrange (),
           .vcounderrange ());
defparam
    altpll_component.clk0_divide_by = 5,
    altpll_component.clk0_duty_cycle = 50,
    altpll_component.clk0_multiply_by = 2,
    altpll_component.clk0_phase_shift = "0",
    altpll_component.compensate_clock = "CLK0",
    altpll_component.inclk0_input_frequency = 10000,
    altpll_component.intended_device_family = "Cyclone II",
    altpll_component.lpm_hint = "CBX_MODULE_PREFIX=pll",
    altpll_component.lpm_type = "altpll",
    altpll_component.operation_mode = "NORMAL",
    altpll_component.port_activeclock = "PORT_UNUSED",
    altpll_component.port_areset = "PORT_UNUSED",
    altpll_component.port_clkbad0 = "PORT_UNUSED",
    altpll_component.port_clkbad1 = "PORT_UNUSED",
    altpll_component.port_clkloss = "PORT_UNUSED",
    altpll_component.port_clkswitch = "PORT_UNUSED",
    altpll_component.port_configupdate = "PORT_UNUSED",
    altpll_component.port_fbin = "PORT_UNUSED",
    altpll_component.port_inclk0 = "PORT_USED",
    altpll_component.port_inclk1 = "PORT_UNUSED",
    altpll_component.port_locked = "PORT_UNUSED",
    altpll_component.port_pfdena = "PORT_UNUSED",
    altpll_component.port_phasecounterselect = "PORT_UNUSED",
    altpll_component.port_phasedone = "PORT_UNUSED",
    altpll_component.port_phasestep = "PORT_UNUSED",
    altpll_component.port_phaseupdown = "PORT_UNUSED",
    altpll_component.port_pllena = "PORT_UNUSED",
    altpll_component.port_scanaclr = "PORT_UNUSED",
    altpll_component.port_scanclk = "PORT_UNUSED",
    altpll_component.port_scanclkena = "PORT_UNUSED",
    altpll_component.port_scandata = "PORT_UNUSED",
    altpll_component.port_scandataout = "PORT_UNUSED",
    altpll_component.port_scandone = "PORT_UNUSED",
    altpll_component.port_scanread = "PORT_UNUSED",
    altpll_component.port_scanwrite = "PORT_UNUSED",
    altpll_component.port_clk0 = "PORT_USED",
    altpll_component.port_clk1 = "PORT_UNUSED",
    altpll_component.port_clk2 = "PORT_UNUSED",
    altpll_component.port_clk3 = "PORT_UNUSED",
    altpll_component.port_clk4 = "PORT_UNUSED",
    altpll_component.port_clk5 = "PORT_UNUSED",
    altpll_component.port_clkena0 = "PORT_UNUSED",
    altpll_component.port_clkena1 = "PORT_UNUSED",
    altpll_component.port_clkena2 = "PORT_UNUSED",
    altpll_component.port_clkena3 = "PORT_UNUSED",
    altpll_component.port_clkena4 = "PORT_UNUSED",
    altpll_component.port_clkena5 = "PORT_UNUSED",
    altpll_component.port_extclk0 = "PORT_UNUSED",
    altpll_component.port_extclk1 = "PORT_UNUSED",
    altpll_component.port_extclk2 = "PORT_UNUSED",
    altpll_component.port_extclk3 = "PORT_UNUSED";


endmodule

    // ============================================================
    // CNX file retrieval info
    // ============================================================
    // Retrieval info: PRIVATE: ACTIVECLK_CHECK STRING "0"
    // Retrieval info: PRIVATE: BANDWIDTH STRING "1.000"
    // Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED STRING "0"
    // Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT STRING "MHz"
    // Retrieval info: PRIVATE: BANDWIDTH_PRESET STRING "Low"
    // Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO STRING "1"
    // Retrieval info: PRIVATE: BANDWIDTH_USE_CUSTOM STRING "0"
    // Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET STRING "0"
    // Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK STRING "0"
    // Retrieval info: PRIVATE: CLKLOSS_CHECK STRING "0"
    // Retrieval info: PRIVATE: CLKSWITCH_CHECK STRING "1"
    // Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO STRING "0"
    // Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK STRING "0"
    // Retrieval info: PRIVATE: CREATE_INCLK1_CHECK STRING "0"
    // Retrieval info: PRIVATE: CUR_DEDICATED_CLK STRING "c0"
    // Retrieval info: PRIVATE: CUR_FBIN_CLK STRING "c0"
    // Retrieval info: PRIVATE: DEVICE_SPEED_GRADE STRING "8"
    // Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "5"
    // Retrieval info: PRIVATE: DUTY_CYCLE0 STRING "50.00000000"
    // Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE0 STRING "40.000000"
    // Retrieval info: PRIVATE: EXPLICIT_SWITCHOVER_COUNTER STRING "0"
    // Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO STRING "0"
    // Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED STRING "1"
    // Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED STRING "1"
    // Retrieval info: PRIVATE: GLOCKED_MODE_CHECK STRING "0"
    // Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "1048575"
    // Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER STRING "1"
    // Retrieval info: PRIVATE: INCLK0_FREQ_EDIT STRING "100.000"
    // Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO STRING "MHz"
    // Retrieval info: PRIVATE: INCLK1_FREQ_EDIT STRING "100.000"
    // Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED STRING "1"
    // Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED STRING "1"
    // Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO STRING "MHz"
    // Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
    // Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO STRING "1"
    // Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK STRING "0"
    // Retrieval info: PRIVATE: LONG_SCAN_RADIO STRING "1"
    // Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE STRING "Not Available"
    // Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
    // Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 STRING "deg"
    // Retrieval info: PRIVATE: MIG_DEVICE_SPEED_GRADE STRING "Any"
    // Retrieval info: PRIVATE: MIRROR_CLK0 STRING "0"
    // Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "2"
    // Retrieval info: PRIVATE: NORMAL_MODE_RADIO STRING "1"
    // Retrieval info: PRIVATE: OUTPUT_FREQ0 STRING "100.00000000"
    // Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 STRING "0"
    // Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 STRING "MHz"
    // Retrieval info: PRIVATE: PHASE_RECONFIG_FEATURE_ENABLED STRING "0"
    // Retrieval info: PRIVATE: PHASE_RECONFIG_INPUTS_CHECK STRING "0"
    // Retrieval info: PRIVATE: PHASE_SHIFT0 STRING "0.00000000"
    // Retrieval info: PRIVATE: PHASE_SHIFT_STEP_ENABLED_CHECK STRING "0"
    // Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 STRING "deg"
    // Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK STRING "0"
    // Retrieval info: PRIVATE: PLL_ARESET_CHECK STRING "0"
    // Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "1"
    // Retrieval info: PRIVATE: PLL_ENA_CHECK STRING "0"
    // Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "0"
    // Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
    // Retrieval info: PRIVATE: PLL_FBMIMIC_CHECK STRING "0"
    // Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
    // Retrieval info: PRIVATE: PLL_PFDENA_CHECK STRING "0"
    // Retrieval info: PRIVATE: PLL_TARGET_HARCOPY_CHECK NUMERIC "0"
    // Retrieval info: PRIVATE: PRIMARY_CLK_COMBO STRING "inclk0"
    // Retrieval info: PRIVATE: RECONFIG_FILE STRING "pll.mif"
    // Retrieval info: PRIVATE: SACN_INPUTS_CHECK STRING "0"
    // Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED STRING "0"
    // Retrieval info: PRIVATE: SELF_RESET_LOCK_LOSS STRING "0"
    // Retrieval info: PRIVATE: SHORT_SCAN_RADIO STRING "0"
    // Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED STRING "0"
    // Retrieval info: PRIVATE: SPREAD_FREQ STRING "50.000"
    // Retrieval info: PRIVATE: SPREAD_FREQ_UNIT STRING "KHz"
    // Retrieval info: PRIVATE: SPREAD_PERCENT STRING "0.500"
    // Retrieval info: PRIVATE: SPREAD_USE STRING "0"
    // Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO STRING "0"
    // Retrieval info: PRIVATE: STICKY_CLK0 STRING "1"
    // Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
    // Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED STRING "1"
    // Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
    // Retrieval info: PRIVATE: USE_CLK0 STRING "1"
    // Retrieval info: PRIVATE: USE_CLKENA0 STRING "0"
    // Retrieval info: PRIVATE: USE_MIL_SPEED_GRADE NUMERIC "0"
    // Retrieval info: PRIVATE: ZERO_DELAY_RADIO STRING "0"
    // Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
    // Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "5"
    // Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
    // Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "2"
    // Retrieval info: CONSTANT: CLK0_PHASE_SHIFT STRING "0"
    // Retrieval info: CONSTANT: COMPENSATE_CLOCK STRING "CLK0"
    // Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "10000"
    // Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
    // Retrieval info: CONSTANT: LPM_TYPE STRING "altpll"
    // Retrieval info: CONSTANT: OPERATION_MODE STRING "NORMAL"
    // Retrieval info: CONSTANT: PORT_ACTIVECLOCK STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_ARESET STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_CLKBAD0 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_CLKBAD1 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_CLKLOSS STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_CLKSWITCH STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_CONFIGUPDATE STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_FBIN STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_INCLK0 STRING "PORT_USED"
    // Retrieval info: CONSTANT: PORT_INCLK1 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_LOCKED STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PFDENA STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PHASECOUNTERSELECT STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PHASEDONE STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PHASESTEP STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PHASEUPDOWN STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_PLLENA STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANACLR STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANCLK STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANCLKENA STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANDATA STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANDATAOUT STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANDONE STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANREAD STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_SCANWRITE STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clk0 STRING "PORT_USED"
    // Retrieval info: CONSTANT: PORT_clk1 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clk2 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clk3 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clk4 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clk5 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena0 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena1 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena2 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena3 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena4 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_clkena5 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_extclk0 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_extclk1 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_extclk2 STRING "PORT_UNUSED"
    // Retrieval info: CONSTANT: PORT_extclk3 STRING "PORT_UNUSED"
    // Retrieval info: USED_PORT: @clk 0 0 6 0 OUTPUT_CLK_EXT VCC "@clk[5..0]"
    // Retrieval info: USED_PORT: @extclk 0 0 4 0 OUTPUT_CLK_EXT VCC "@extclk[3..0]"
    // Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT_CLK_EXT VCC "c0"
    // Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT_CLK_EXT GND "inclk0"
    // Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
    // Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
    // Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll.v TRUE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll.ppf TRUE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll.inc FALSE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll.cmp FALSE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll.bsf FALSE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll_inst.v FALSE
    // Retrieval info: GEN_FILE: TYPE_NORMAL pll_bb.v FALSE
    // Retrieval info: LIB_FILE: altera_mf
    // Retrieval info: CBX_MODULE_PREFIX: ON
